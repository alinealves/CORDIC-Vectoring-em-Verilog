library verilog;
use verilog.vl_types.all;
entity AJ_vlg_vec_tst is
end AJ_vlg_vec_tst;
